`include "definitions.vh"
module iExecute_test;
reg [`WORD-1:0] pc_in, read_data1, read_data2, sign_extend;
reg [10:0] opcode;
reg [1:0] alu_op;
reg alu_src;
wire [`WORD-1:0] alu_result, branch_target;
wire zero;


endmodule